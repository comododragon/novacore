// NovaCOREBlaster.v

// Generated using ACDS version 14.1 186 at 2017.03.31.13:08:48

`timescale 1 ps / 1 ps
module NovaCOREBlaster (
		output wire [27:0] c_bus_export,       //       c_bus.export
		output wire        c_clk_export,       //       c_clk.export
		output wire [3:0]  c_dimension_export, // c_dimension.export
		output wire        c_dimswitch_export, // c_dimswitch.export
		output wire [3:0]  c_uid_export,       //       c_uid.export
		input  wire        clk_clk,            //         clk.clk
		output wire        mode_export,        //        mode.export
		input  wire        reset_reset_n       //       reset.reset_n
	);

	wire  [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [20:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [20:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_pio_mode_s1_chipselect;                  // mm_interconnect_0:pio_mode_s1_chipselect -> pio_mode:chipselect
	wire  [31:0] mm_interconnect_0_pio_mode_s1_readdata;                    // pio_mode:readdata -> mm_interconnect_0:pio_mode_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_mode_s1_address;                     // mm_interconnect_0:pio_mode_s1_address -> pio_mode:address
	wire         mm_interconnect_0_pio_mode_s1_write;                       // mm_interconnect_0:pio_mode_s1_write -> pio_mode:write_n
	wire  [31:0] mm_interconnect_0_pio_mode_s1_writedata;                   // mm_interconnect_0:pio_mode_s1_writedata -> pio_mode:writedata
	wire         mm_interconnect_0_pio_c_bus_s1_chipselect;                 // mm_interconnect_0:pio_c_bus_s1_chipselect -> pio_c_bus:chipselect
	wire  [31:0] mm_interconnect_0_pio_c_bus_s1_readdata;                   // pio_c_bus:readdata -> mm_interconnect_0:pio_c_bus_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_c_bus_s1_address;                    // mm_interconnect_0:pio_c_bus_s1_address -> pio_c_bus:address
	wire         mm_interconnect_0_pio_c_bus_s1_write;                      // mm_interconnect_0:pio_c_bus_s1_write -> pio_c_bus:write_n
	wire  [31:0] mm_interconnect_0_pio_c_bus_s1_writedata;                  // mm_interconnect_0:pio_c_bus_s1_writedata -> pio_c_bus:writedata
	wire         mm_interconnect_0_pio_c_dimswitch_s1_chipselect;           // mm_interconnect_0:pio_c_dimswitch_s1_chipselect -> pio_c_dimswitch:chipselect
	wire  [31:0] mm_interconnect_0_pio_c_dimswitch_s1_readdata;             // pio_c_dimswitch:readdata -> mm_interconnect_0:pio_c_dimswitch_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_c_dimswitch_s1_address;              // mm_interconnect_0:pio_c_dimswitch_s1_address -> pio_c_dimswitch:address
	wire         mm_interconnect_0_pio_c_dimswitch_s1_write;                // mm_interconnect_0:pio_c_dimswitch_s1_write -> pio_c_dimswitch:write_n
	wire  [31:0] mm_interconnect_0_pio_c_dimswitch_s1_writedata;            // mm_interconnect_0:pio_c_dimswitch_s1_writedata -> pio_c_dimswitch:writedata
	wire         mm_interconnect_0_pio_c_dimension_s1_chipselect;           // mm_interconnect_0:pio_c_dimension_s1_chipselect -> pio_c_dimension:chipselect
	wire  [31:0] mm_interconnect_0_pio_c_dimension_s1_readdata;             // pio_c_dimension:readdata -> mm_interconnect_0:pio_c_dimension_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_c_dimension_s1_address;              // mm_interconnect_0:pio_c_dimension_s1_address -> pio_c_dimension:address
	wire         mm_interconnect_0_pio_c_dimension_s1_write;                // mm_interconnect_0:pio_c_dimension_s1_write -> pio_c_dimension:write_n
	wire  [31:0] mm_interconnect_0_pio_c_dimension_s1_writedata;            // mm_interconnect_0:pio_c_dimension_s1_writedata -> pio_c_dimension:writedata
	wire         mm_interconnect_0_bitstream_memory_s1_chipselect;          // mm_interconnect_0:bitstream_memory_s1_chipselect -> bitstream_memory:chipselect
	wire  [31:0] mm_interconnect_0_bitstream_memory_s1_readdata;            // bitstream_memory:readdata -> mm_interconnect_0:bitstream_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_bitstream_memory_s1_address;             // mm_interconnect_0:bitstream_memory_s1_address -> bitstream_memory:address
	wire   [3:0] mm_interconnect_0_bitstream_memory_s1_byteenable;          // mm_interconnect_0:bitstream_memory_s1_byteenable -> bitstream_memory:byteenable
	wire         mm_interconnect_0_bitstream_memory_s1_write;               // mm_interconnect_0:bitstream_memory_s1_write -> bitstream_memory:write
	wire  [31:0] mm_interconnect_0_bitstream_memory_s1_writedata;           // mm_interconnect_0:bitstream_memory_s1_writedata -> bitstream_memory:writedata
	wire         mm_interconnect_0_bitstream_memory_s1_clken;               // mm_interconnect_0:bitstream_memory_s1_clken -> bitstream_memory:clken
	wire         mm_interconnect_0_pio_c_clk_s1_chipselect;                 // mm_interconnect_0:pio_c_clk_s1_chipselect -> pio_c_clk:chipselect
	wire  [31:0] mm_interconnect_0_pio_c_clk_s1_readdata;                   // pio_c_clk:readdata -> mm_interconnect_0:pio_c_clk_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_c_clk_s1_address;                    // mm_interconnect_0:pio_c_clk_s1_address -> pio_c_clk:address
	wire         mm_interconnect_0_pio_c_clk_s1_write;                      // mm_interconnect_0:pio_c_clk_s1_write -> pio_c_clk:write_n
	wire  [31:0] mm_interconnect_0_pio_c_clk_s1_writedata;                  // mm_interconnect_0:pio_c_clk_s1_writedata -> pio_c_clk:writedata
	wire         mm_interconnect_0_pio_c_uid_s1_chipselect;                 // mm_interconnect_0:pio_c_uid_s1_chipselect -> pio_c_uid:chipselect
	wire  [31:0] mm_interconnect_0_pio_c_uid_s1_readdata;                   // pio_c_uid:readdata -> mm_interconnect_0:pio_c_uid_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_c_uid_s1_address;                    // mm_interconnect_0:pio_c_uid_s1_address -> pio_c_uid:address
	wire         mm_interconnect_0_pio_c_uid_s1_write;                      // mm_interconnect_0:pio_c_uid_s1_write -> pio_c_uid:write_n
	wire  [31:0] mm_interconnect_0_pio_c_uid_s1_writedata;                  // mm_interconnect_0:pio_c_uid_s1_writedata -> pio_c_uid:writedata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [bitstream_memory:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, onchip_memory2:reset, pio_c_bus:reset_n, pio_c_clk:reset_n, pio_c_dimension:reset_n, pio_c_dimswitch:reset_n, pio_c_uid:reset_n, pio_mode:reset_n, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [bitstream_memory:reset_req, nios2_gen2:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> rst_controller:reset_in1

	NovaCOREBlaster_bitstream_memory bitstream_memory (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_bitstream_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_bitstream_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_bitstream_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_bitstream_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_bitstream_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_bitstream_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_bitstream_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	NovaCOREBlaster_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	NovaCOREBlaster_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	NovaCOREBlaster_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)              //       .reset_req
	);

	NovaCOREBlaster_pio_c_bus pio_c_bus (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_c_bus_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_c_bus_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_c_bus_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_c_bus_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_c_bus_s1_readdata),   //                    .readdata
		.out_port   (c_bus_export)                               // external_connection.export
	);

	NovaCOREBlaster_pio_c_clk pio_c_clk (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_c_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_c_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_c_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_c_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_c_clk_s1_readdata),   //                    .readdata
		.out_port   (c_clk_export)                               // external_connection.export
	);

	NovaCOREBlaster_pio_c_dimension pio_c_dimension (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_pio_c_dimension_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_c_dimension_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_c_dimension_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_c_dimension_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_c_dimension_s1_readdata),   //                    .readdata
		.out_port   (c_dimension_export)                               // external_connection.export
	);

	NovaCOREBlaster_pio_c_clk pio_c_dimswitch (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_pio_c_dimswitch_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_c_dimswitch_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_c_dimswitch_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_c_dimswitch_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_c_dimswitch_s1_readdata),   //                    .readdata
		.out_port   (c_dimswitch_export)                               // external_connection.export
	);

	NovaCOREBlaster_pio_c_dimension pio_c_uid (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_c_uid_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_c_uid_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_c_uid_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_c_uid_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_c_uid_s1_readdata),   //                    .readdata
		.out_port   (c_uid_export)                               // external_connection.export
	);

	NovaCOREBlaster_pio_mode pio_mode (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_mode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_mode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_mode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_mode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_mode_s1_readdata),   //                    .readdata
		.out_port   (mode_export)                               // external_connection.export
	);

	NovaCOREBlaster_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	NovaCOREBlaster_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                               (clk_clk),                                                   //                             clk_50_clk.clk
		.nios2_gen2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios2_gen2_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address               (nios2_gen2_data_master_address),                            //                 nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest           (nios2_gen2_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_gen2_data_master_byteenable            (nios2_gen2_data_master_byteenable),                         //                                       .byteenable
		.nios2_gen2_data_master_read                  (nios2_gen2_data_master_read),                               //                                       .read
		.nios2_gen2_data_master_readdata              (nios2_gen2_data_master_readdata),                           //                                       .readdata
		.nios2_gen2_data_master_write                 (nios2_gen2_data_master_write),                              //                                       .write
		.nios2_gen2_data_master_writedata             (nios2_gen2_data_master_writedata),                          //                                       .writedata
		.nios2_gen2_data_master_debugaccess           (nios2_gen2_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_gen2_instruction_master_address        (nios2_gen2_instruction_master_address),                     //          nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest    (nios2_gen2_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_gen2_instruction_master_read           (nios2_gen2_instruction_master_read),                        //                                       .read
		.nios2_gen2_instruction_master_readdata       (nios2_gen2_instruction_master_readdata),                    //                                       .readdata
		.bitstream_memory_s1_address                  (mm_interconnect_0_bitstream_memory_s1_address),             //                    bitstream_memory_s1.address
		.bitstream_memory_s1_write                    (mm_interconnect_0_bitstream_memory_s1_write),               //                                       .write
		.bitstream_memory_s1_readdata                 (mm_interconnect_0_bitstream_memory_s1_readdata),            //                                       .readdata
		.bitstream_memory_s1_writedata                (mm_interconnect_0_bitstream_memory_s1_writedata),           //                                       .writedata
		.bitstream_memory_s1_byteenable               (mm_interconnect_0_bitstream_memory_s1_byteenable),          //                                       .byteenable
		.bitstream_memory_s1_chipselect               (mm_interconnect_0_bitstream_memory_s1_chipselect),          //                                       .chipselect
		.bitstream_memory_s1_clken                    (mm_interconnect_0_bitstream_memory_s1_clken),               //                                       .clken
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.nios2_gen2_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //             nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                       .write
		.nios2_gen2_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                       .read
		.nios2_gen2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_gen2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_gen2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.onchip_memory2_s1_address                    (mm_interconnect_0_onchip_memory2_s1_address),               //                      onchip_memory2_s1.address
		.onchip_memory2_s1_write                      (mm_interconnect_0_onchip_memory2_s1_write),                 //                                       .write
		.onchip_memory2_s1_readdata                   (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                       .readdata
		.onchip_memory2_s1_writedata                  (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                       .writedata
		.onchip_memory2_s1_byteenable                 (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                       .byteenable
		.onchip_memory2_s1_chipselect                 (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                       .chipselect
		.onchip_memory2_s1_clken                      (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                       .clken
		.pio_c_bus_s1_address                         (mm_interconnect_0_pio_c_bus_s1_address),                    //                           pio_c_bus_s1.address
		.pio_c_bus_s1_write                           (mm_interconnect_0_pio_c_bus_s1_write),                      //                                       .write
		.pio_c_bus_s1_readdata                        (mm_interconnect_0_pio_c_bus_s1_readdata),                   //                                       .readdata
		.pio_c_bus_s1_writedata                       (mm_interconnect_0_pio_c_bus_s1_writedata),                  //                                       .writedata
		.pio_c_bus_s1_chipselect                      (mm_interconnect_0_pio_c_bus_s1_chipselect),                 //                                       .chipselect
		.pio_c_clk_s1_address                         (mm_interconnect_0_pio_c_clk_s1_address),                    //                           pio_c_clk_s1.address
		.pio_c_clk_s1_write                           (mm_interconnect_0_pio_c_clk_s1_write),                      //                                       .write
		.pio_c_clk_s1_readdata                        (mm_interconnect_0_pio_c_clk_s1_readdata),                   //                                       .readdata
		.pio_c_clk_s1_writedata                       (mm_interconnect_0_pio_c_clk_s1_writedata),                  //                                       .writedata
		.pio_c_clk_s1_chipselect                      (mm_interconnect_0_pio_c_clk_s1_chipselect),                 //                                       .chipselect
		.pio_c_dimension_s1_address                   (mm_interconnect_0_pio_c_dimension_s1_address),              //                     pio_c_dimension_s1.address
		.pio_c_dimension_s1_write                     (mm_interconnect_0_pio_c_dimension_s1_write),                //                                       .write
		.pio_c_dimension_s1_readdata                  (mm_interconnect_0_pio_c_dimension_s1_readdata),             //                                       .readdata
		.pio_c_dimension_s1_writedata                 (mm_interconnect_0_pio_c_dimension_s1_writedata),            //                                       .writedata
		.pio_c_dimension_s1_chipselect                (mm_interconnect_0_pio_c_dimension_s1_chipselect),           //                                       .chipselect
		.pio_c_dimswitch_s1_address                   (mm_interconnect_0_pio_c_dimswitch_s1_address),              //                     pio_c_dimswitch_s1.address
		.pio_c_dimswitch_s1_write                     (mm_interconnect_0_pio_c_dimswitch_s1_write),                //                                       .write
		.pio_c_dimswitch_s1_readdata                  (mm_interconnect_0_pio_c_dimswitch_s1_readdata),             //                                       .readdata
		.pio_c_dimswitch_s1_writedata                 (mm_interconnect_0_pio_c_dimswitch_s1_writedata),            //                                       .writedata
		.pio_c_dimswitch_s1_chipselect                (mm_interconnect_0_pio_c_dimswitch_s1_chipselect),           //                                       .chipselect
		.pio_c_uid_s1_address                         (mm_interconnect_0_pio_c_uid_s1_address),                    //                           pio_c_uid_s1.address
		.pio_c_uid_s1_write                           (mm_interconnect_0_pio_c_uid_s1_write),                      //                                       .write
		.pio_c_uid_s1_readdata                        (mm_interconnect_0_pio_c_uid_s1_readdata),                   //                                       .readdata
		.pio_c_uid_s1_writedata                       (mm_interconnect_0_pio_c_uid_s1_writedata),                  //                                       .writedata
		.pio_c_uid_s1_chipselect                      (mm_interconnect_0_pio_c_uid_s1_chipselect),                 //                                       .chipselect
		.pio_mode_s1_address                          (mm_interconnect_0_pio_mode_s1_address),                     //                            pio_mode_s1.address
		.pio_mode_s1_write                            (mm_interconnect_0_pio_mode_s1_write),                       //                                       .write
		.pio_mode_s1_readdata                         (mm_interconnect_0_pio_mode_s1_readdata),                    //                                       .readdata
		.pio_mode_s1_writedata                        (mm_interconnect_0_pio_mode_s1_writedata),                   //                                       .writedata
		.pio_mode_s1_chipselect                       (mm_interconnect_0_pio_mode_s1_chipselect),                  //                                       .chipselect
		.timer_s1_address                             (mm_interconnect_0_timer_s1_address),                        //                               timer_s1.address
		.timer_s1_write                               (mm_interconnect_0_timer_s1_write),                          //                                       .write
		.timer_s1_readdata                            (mm_interconnect_0_timer_s1_readdata),                       //                                       .readdata
		.timer_s1_writedata                           (mm_interconnect_0_timer_s1_writedata),                      //                                       .writedata
		.timer_s1_chipselect                          (mm_interconnect_0_timer_s1_chipselect)                      //                                       .chipselect
	);

	NovaCOREBlaster_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
